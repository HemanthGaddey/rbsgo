module ir_test(
	input clk_50_,
	input dout_,
	output adc_cs_n_,
	output din_,
	output adc_sck_,
	
	output led1_,
	output led2_,
	output led3_,
	output led4_,
	output led5_,
	output led6_,
	output led7_,
	output led8_
	);
	
	reg led1,led2,led3,led4,led5,led6,led7,led8;
	wire [11:0]ir1;
	wire [11:0]ir2;
	wire [11:0]ir3;
	assign led1_ = led1;
	assign led2_ = led2;
	assign led3_ = led3;
	assign led4_ = led4;
	assign led5_ = led5;
	assign led6_ = led6;
	assign led7_ = led7;
	assign led8_ = led8;
	
	adc_control ac(
		.clk_50(clk_50_),
		.dout(dout_),
		.adc_cs_n(adc_cs_n_),
		.din(din_),
		.adc_sck(adc_sck_),
		.d_out_ch5(ir1),
		.d_out_ch6(ir2),
		.d_out_ch7(ir3)
	);
	
	
	always @ (posedge clk_50_)	begin
		led1 <= ir1[0];
		led2 <= ir1[1];
		led3 <= ir1[2];
		led4 <= ir1[3];
		led5 <= ir1[4];
		led6 <= ir1[5];
		led7 <= ir1[6];
		led8 <= ir1[7];
	end
	
	endmodule