module motor_test(
	input clk,
	output a1,
	output a2,
	output b1,
	output b2
	);
	assign b1 = 1;
	assign b2 = 0;
	assign a1 = 1;
	assign a2 = 0;
	
	endmodule